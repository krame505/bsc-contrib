package SizedVector where

-- TODO: Where should this library live?
-- It is used in both the COBS and GenC libraries, which are otherwise independent.

import Vector
import Array

type SizeBits n = TLog (TAdd 1 n)

-- Represents a variable-sized vector of max length n
struct SizedVector n a = 
  size :: UInt (SizeBits n)
  items :: Vector n a
 deriving (Eq, Bits)

nil :: SizedVector n a
nil = SizedVector { size=0; items=replicate _; }

fromFullVector :: Vector n a -> SizedVector n a
fromFullVector v = SizedVector { size=fromInteger $ valueOf n; items=v; }

class AppendSizedVector n1 n2 n | n1 n2 -> n where
  append :: SizedVector n1 a -> SizedVector n2 a -> SizedVector n a

instance (Add n1 n2 n, 
          Add p1 (SizeBits n1) (SizeBits n), 
          Add p2 (SizeBits n2) (SizeBits n)) =>
         AppendSizedVector n1 n2 n where
    append :: SizedVector n1 a -> SizedVector n2 a -> SizedVector n a
    append v1 v2 = SizedVector {
      size = zeroExtend v1.size + zeroExtend v2.size;
      items = foldr
        (\ (i, x) result -> update result ((zeroExtend v1.size + fromInteger i) :: UInt (SizeBits n)) x)
        (Vector.append v1.items newVector)
        (zip genVector v2.items);
    }

class ConcatSizedVector n1 n2 n | n1 n2 -> n where
  concat :: Vector n1 (SizedVector n2 a) -> SizedVector n a

instance ConcatSizedVector 0 n 0 where
  concat _ = nil

instance (ConcatSizedVector n1' n2 n', Add n1' 1 n1, AppendSizedVector n' n2 n) =>
         ConcatSizedVector n1 n2 n where
  concat v = append (concat $ init v) $ last v

extend :: (AppendSizedVector n k m) => SizedVector n a -> SizedVector m a
extend v = SizedVector { size = zeroExtend v.size; items = Vector.append v.items $ replicate _; }

accum :: (Add n k m) => Vector n a -> SizedVector m a -> SizedVector m a
accum items v = SizedVector {
  size = v.size + fromInteger (valueOf n);
  items = foldr
    (\ (i, x) result -> update result (v.size + fromInteger i) x)
    v.items (zip genVector items);
}