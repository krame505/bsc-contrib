package SizedVector where

-- TODO: Where should this library live?
-- It is used in both the COBS and GenC libraries, which are otherwise independent.

import Vector

type SizeBits n = TLog (TAdd 1 n)

-- Represents a variable-sized vector of max length n
struct SizedVector n a = 
  size :: UInt (SizeBits n)
  items :: Vector n a
 deriving (Eq, Bits)

nil :: SizedVector n a
nil = SizedVector { size=0; items=replicate _; }

fromFullVector :: Vector n a -> SizedVector n a
fromFullVector v = SizedVector { size=fromInteger $ valueOf n; items=v; }

class AppendSizedVector n1 n2 n | n1 n2 -> n where
  append :: SizedVector n1 a -> SizedVector n2 a -> SizedVector n a

instance (Add n1 n2 n, 
          Add p1 (TLog (TAdd 1 n1)) (SizeBits n), 
          Add p2 (TLog (TAdd 1 n2)) (SizeBits n)) =>
         AppendSizedVector n1 n2 n where
    append :: SizedVector n1 a -> SizedVector n2 a -> SizedVector n a
    append v1 v2 = SizedVector {
      size = zeroExtend v1.size + zeroExtend v2.size;
      items =
        let options :: Vector (TAdd 1 n1) (Vector n a) =
              genWith $ \ i ->
                genWith $ \ j ->
                  if j < i
                  then v1.items !! j
                  else if j < i + valueOf n2
                  then v2.items !! (j - i)
                  else _;
        in select options v1.size;
    }

class ConcatSizedVector n m o | n m -> o where
  concat :: Vector n (SizedVector m a) -> SizedVector o a

instance ConcatSizedVector 0 m 0 where
  concat _ = nil

instance ConcatSizedVector 1 m m where
  concat v = head v

instance (Div n 2 n1, Add n1 n2 n,
          ConcatSizedVector n1 m o1, ConcatSizedVector n2 m o2, AppendSizedVector o1 o2 o) =>
         ConcatSizedVector n m o where
  concat :: Vector n (SizedVector m a) -> SizedVector o a
  concat v =
    let v1 :: Vector n1 (SizedVector m a) = take v
        v2 :: Vector n2 (SizedVector m a) = drop v
    in append (concat v1) (concat v2)

extend :: (AppendSizedVector n k m) => SizedVector n a -> SizedVector m a
extend v = append v $ fromFullVector $ replicate _
